LIBRARY ieee;
USE ieee.std_logic_1164.all; 

ENTITY Tarea2 IS PORT (
	SW  : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
   KEY : IN STD_LOGIC_VECTOR (3 DOWNTO 0);	
	LEDG: OUT STD_LOGIC_VECTOR(0 DOWNTO 0)
);
END Tarea2;

ARCHITECTURE Mux4_1 OF Tarea2 IS
BEGIN
	WITH SW SELECT 
		LEDG(0) <=	NOT KEY(0) WHEN "00",
						NOT KEY(1) WHEN "01",
						NOT KEY(2) WHEN "10",
						NOT KEY(3) WHEN "11";
   
END Mux4_1;